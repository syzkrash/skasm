// Generated with gen_op.vsh on 3rd Jun 2022 18:14:13 (+2)
module assembler
const opmap = {
	"NOOP": u8(0),
	"PANIC": u8(1),
	"DROP": u8(16),
	"DUP": u8(20),
	"SWAP": u8(17),
	"ROT": u8(18),
	"OVER": u8(19),
	"PUSHB": u8(26),
	"PUSHP": u8(27),
	"PUSHI": u8(28),
	"PUSHF": u8(29),
	"PUSHL": u8(30),
	"GETB": u8(32),
	"SETB": u8(33),
	"GETP": u8(34),
	"SETP": u8(35),
	"GETI": u8(36),
	"SETI": u8(37),
	"GETF": u8(38),
	"SETF": u8(39),
	"ADD": u8(48),
	"SUB": u8(49),
	"MUL": u8(50),
	"DIMD": u8(51),
	"LSH": u8(52),
	"RSH": u8(53),
	"AND": u8(54),
	"OR": u8(55),
	"XOR": u8(56),
	"NOT": u8(57),
	"LABEL": u8(64),
	"FUNC": u8(65),
	"JMP": u8(66),
	"CALL": u8(67),
	"RET": u8(68),
	"JMPIF": u8(79),
}
